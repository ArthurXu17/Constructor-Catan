RED
0 1 1 1 1 r h 30 H 20 H 
1 1 2 1 1 r h 13 B 53 B 
1 0 2 1 1 r h 25 T 23 B 5 B 
1 0 1 0 0 r h 49 B 35 B 
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9 
13