RED
0 0 0 0 1 r h 45 B 5 B 
0 1 1 0 1 r h 40 B 15 B 
0 0 0 0 0 r h 35 B 20 B 
0 0 2 1 0 r h 30 B 25 B 
0 2 0 3 0 3 0 4 1 4 1 5 1 5 1 6 2 6 5 7 2 8 2 8 2 9 3 9 3 10 3 10 4 11 4 11 4 12 
9