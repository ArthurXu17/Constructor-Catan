BLUE
1 0 0 0 0 r h 20 B 0 B 
0 0 0 0 0 r h 18 B 2 B 
1 0 0 0 0 r h 15 B 5 B 
1 0 0 0 0 r h 11 B 8 B 
3 5 4 6 1 8 2 10 0 4 2 5 2 2 1 3 2 11 3 8 4 12 4 10 1 9 0 4 5 7 3 9 0 3 0 6 1 11 
14