BLUE
1 1 1 1 0 r 21 18 h 19 B 32 B 
1 1 4 2 2 r 68 h 50 B 52 B 
2 1 2 3 1 r h 44 B 48 H 
10 10 10 10 10 r h 0 B 4 H 
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9 
4