BLUE
0 0 0 0 0 r h 
0 0 0 0 0 r h 
0 0 0 0 0 r h 
0 0 0 0 0 r h 
3 10 4 8 5 7 4 3 2 6 0 6 1 11 0 10 2 11 2 9 0 4 1 12 4 8 1 5 3 3 3 9 2 5 0 2 1 4 
2