RED
6 0 0 0 0 r h 51 B 40 B 8 H 4 T 52 B 0 B 
0 0 3 0 1 r 56 h 44 B 13 T 
0 0 0 0 0 r h 30 B 
0 3 1 0 0 r h 25 T 2 H 
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9 
8