BLUE
499 514 521 496 533 r h 36 T 24 H 12 B 
499 514 521 496 533 r h 31 T 19 H 7 B 
533 501 493 493 544 r 49 57 h 33 T 21 H 9 B 
535 502 492 494 542 r h 35 T 23 H 11 B 
0 3 1 10 3 5 1 4 5 7 3 10 2 11 0 3 3 8 0 2 0 6 1 8 4 12 1 5 4 11 2 4 4 6 2 9 2 9 
4